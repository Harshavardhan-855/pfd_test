magic
tech sky130A
timestamp 1708506111
<< checkpaint >>
rect -630 -330 2215 2037
rect -630 -1630 730 -330
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
rect 0 -600 100 -500
rect 0 -800 100 -700
rect 0 -1000 100 -900
use pfd  x1
timestamp 1708506044
transform 1 0 -393 0 1 1240
box 393 -940 1978 167
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 128 0 0 0 A1
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 128 0 0 0 B1
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 128 0 0 0 QA1
port 2 nsew
flabel metal1 0 -600 100 -500 0 FreeSans 128 0 0 0 QB1
port 3 nsew
flabel metal1 0 -800 100 -700 0 FreeSans 128 0 0 0 VDD1
port 4 nsew
flabel metal1 0 -1000 100 -900 0 FreeSans 128 0 0 0 VSS1
port 5 nsew
<< end >>
